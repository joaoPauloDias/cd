library verilog;
use verilog.vl_types.all;
entity jpd_generic_ula_vlg_vec_tst is
end jpd_generic_ula_vlg_vec_tst;
