library verilog;
use verilog.vl_types.all;
entity jpd_mux_2x1_8bit_vlg_vec_tst is
end jpd_mux_2x1_8bit_vlg_vec_tst;
