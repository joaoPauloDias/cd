library verilog;
use verilog.vl_types.all;
entity jpd_counter_8_vlg_vec_tst is
end jpd_counter_8_vlg_vec_tst;
