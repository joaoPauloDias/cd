library verilog;
use verilog.vl_types.all;
entity jpd_s8bit_vlg_check_tst is
    port(
        co              : in     vl_logic;
        s               : in     vl_logic_vector(7 downto 0);
        sampler_rx      : in     vl_logic
    );
end jpd_s8bit_vlg_check_tst;
