library verilog;
use verilog.vl_types.all;
entity jpd_mux_4x1_vlg_check_tst is
    port(
        s               : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end jpd_mux_4x1_vlg_check_tst;
