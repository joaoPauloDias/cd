library verilog;
use verilog.vl_types.all;
entity jpd_mux_8x1_vlg_vec_tst is
end jpd_mux_8x1_vlg_vec_tst;
