library verilog;
use verilog.vl_types.all;
entity jpd_control_vlg_vec_tst is
end jpd_control_vlg_vec_tst;
