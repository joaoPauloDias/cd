library verilog;
use verilog.vl_types.all;
entity jpd_counter_display_vlg_vec_tst is
end jpd_counter_display_vlg_vec_tst;
