library verilog;
use verilog.vl_types.all;
entity jpd_fsm_vlg_vec_tst is
end jpd_fsm_vlg_vec_tst;
