library verilog;
use verilog.vl_types.all;
entity jpd_mux_4x1_vlg_vec_tst is
end jpd_mux_4x1_vlg_vec_tst;
