library verilog;
use verilog.vl_types.all;
entity jpd_ha_vlg_vec_tst is
end jpd_ha_vlg_vec_tst;
