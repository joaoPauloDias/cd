library verilog;
use verilog.vl_types.all;
entity jpd_neg_8bit_vlg_vec_tst is
end jpd_neg_8bit_vlg_vec_tst;
