library verilog;
use verilog.vl_types.all;
entity jpd_fa_vlg_vec_tst is
end jpd_fa_vlg_vec_tst;
