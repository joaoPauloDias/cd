library verilog;
use verilog.vl_types.all;
entity jpd_neg_8bit_vlg_sample_tst is
    port(
        A               : in     vl_logic_vector(7 downto 0);
        sampler_tx      : out    vl_logic
    );
end jpd_neg_8bit_vlg_sample_tst;
