library verilog;
use verilog.vl_types.all;
entity jpd_s8bit_vlg_vec_tst is
end jpd_s8bit_vlg_vec_tst;
